
----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:31:53 11/28/2017 
-- Design Name: 
-- Module Name:    InstructionMemory - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity InstructionMemory is
port(
     skey: in std_logic_vector(127 downto 0);
	  din: in std_logic_vector(63 downto 0);
     address: in std_logic_vector(31 downto 0);
	 mode: in std_logic;
	  Instruction: out std_logic_vector(31 downto 0);
	  	 ins_num: out integer);
	  
end InstructionMemory;

architecture Behavioral of InstructionMemory is

type ramtype3 is array(0 to 1056)of std_logic_vector(31 downto 0);
signal imem: ramtype3:=
(
"00000000000000000000100000010000",--0 ADD RO,RO, R1 R1=0
"00000000000000000001000000010000",--1 ADD R0,RO, R2 R2=0
"00000000000000000001100000010000",--2 ADD RO,RO, R3 R3=0
"00000100000111100000000000000000",--3 ****ADDI,RO,R30,skey(31 downto 16) R30=XXX..skey(31 downto 16)
"00010111110111100000000000010000",--4 SHL R30 R30 16 R30=skey(31 downto 16)...000
"00000100000111010000000000000000",--5 ****ADDI,RO,R29,SKEY(15 downto 0) R29=XXX��..skey(15 downto 0)
"00010111101111010000000000010000",--6 SHL R29 R29 16 R29=skey(15 downto 0)��000     remove sign extension
"00011011101111010000000000010000",--7 SHR R29 R29 16 R29=000��..skey(15 downto 0)     remove sign extension
"00000011110111011111000000010000",--8 ADD,R30 R29,R30 R30=skey(31 downto 0) 
"00100000000111100000000000011010",--9 SW RO, R30 offset M[0+offset1]<-R30
"00000100000111100000000000000000",--10 *****ADDI,RO,R30,skey(63 downto 48) R30=XXX..skey(63 downto 48)
"00010111110111100000000000010000",--11 SHL R30 R30 16 R30=skey(63 downto 48)...000
"00000100000111010000000000000000",--12 **** ADDI,RO,R29,SKEY(47 downto 32) R29=XXX��..skey(47 downto 32)
"00010111101111010000000000010000",--13 SHL R29 R29 16 R29=skey(47 downto 32)��000     remove sign extension
"00011011101111010000000000010000",--14 SHR R29 R29 16 R29=000��..skey(47 downto 32)     remove sign extension
"00000011110111011111000000010000",--15 ADD,R30 R29,R30 R30=skey(63 downto 32) 
"00100000000111100000000000011011",--16 SW RO, R30 offset M[0+offset2]<-R30
"00000100000111100000000000000000",--17 ****ADDI,RO,R30,skey(95 downto 80) R30=XXX..skey(95 downto 80)
"00010111110111100000000000010000",--18 SHL R30 R30 16 R30=skey(95 downto 80)...000
"00000100000111010000000000000000",--19 **** ADDI,RO,R29,SKEY(79 downto 64) R29=XXX��..skey(79 downto 64)
"00010111101111010000000000010000",--20 SHL R29 R29 16 R29=skey(79 downto 64)��000     remove sign extension
"00011011101111010000000000010000",--21 SHR R29 R29 16 R29=000��..skey(79 downto 64)     remove sign extension
"00000011110111011111000000010000",--22 ADD,R30 R29,R30 R30=skey(95 downto 64) 
"00100000000111100000000000011100",--23 SW RO, R30 offset M[0+offset3]<-R30
"00000100000111100000000000000000",--24 ******ADDI,RO,R30,skey(127 downto 112) R30=XXX..skey(127 downto 112)
"00010111110111100000000000010000",--25 SHL R30 R30 16 R30=skey(127 downto 112)...000
"00000100000111010000000000000000",--26******* ADDI,RO,R29,SKEY(111 downto 96) R29=XXX��..skey(111 downto 96)
"00010111101111010000000000010000",--27 SHL R29 R29 16 R29=skey(111 downto 96)��000     remove sign extension
"00011011101111010000000000010000",--28 SHR R29 R29 16 R29=000��..skey(111 downto 96)     remove sign extension
"00000011110111011111000000010000",--29 ADD,R30 R29,R30 R30=skey(127 downto 96) 
"00100000000111100000000000011101",--30 SW RO, R30 offset M[0+offset4]<-R30
"00000100000101010000000000000100",--31 ADDI,RO,R21,4 R21=4
"00000100000101100000000000011010",--32 ADDI RO R22,26 R22=26
"00000100000101110000000001001110",--33 ADDI R0 R23,78 R23=78
"00000000000000000010000000010000",--34 ADD RO RO R4 R4=0
"00000000000000000010100000010000",--35 ADD RO RO R5 R5=0
"00011100010010000000000000000000",--36 R8<-MEM[R2+IMM_S) S[i]
"00011100001010010000000000011010",--37 R9<-MEM(R1+IMM_l) L[j]
"00000000100001010011000000010000",--38 ADD R4 R5,R6  A+B
"00000001000001100101000000010000",--39 ADD R8 R6 R10 A+B+S[i]
																												--"00000100000010110000000000000011",--40 ADDI RO R11 3 
"00000000000000000110000000010000",--40 ADD RO RO R12
																												--"00101001011011000000000000000101",--42 BEQ R11 R12 IMM go to 48
"00010101010011010000000000000011",--41 SHL R10 R13 3
"00011001010011100000000000011101",--42 SHR R10 R14 29
"00000001101011100101000000010000",--43 ADD R13 R14 R10  rotate 1 bit of R10, do it 3 times 	
																												--"00000101100011000000000000000001",--46 ADDI R12 R12 1
																												--"00110000000000000000000000101010",--47 JMP IMM go to 42
"00100000010010100000000000000000",--44 SW R2 R10 IMM_S branch here update S[i]
"00000000000010100010000000010000",--45 add RO R10 R4 put value of A into R4
"00000000100001010011000000010000",--46 add R4 R5 R6 A + B
"00000001001001100101000000010000",--47 add R9 R6 R10 R10 = L[i] + A + B
"00001100110010110000000000011111",--48 ANDI R6 R11 00....11111

																												--"00000000000000000110000000010000",--53 AND RO RO R12
																												--"00101001011011000000000000000101",--54 bEQ R11 R12 IMM
																												--"00010101010011010000000000000001",--55 SHL R10 R13 1
																												--"00011001010011100000000000011111",--56 SHR R10 R14 31
																												--"00000001101011100101000000010000",--57 ADD R13 R14 R10
																												--"00000101100011000000000000000001",--58 ADDI R12 R12 1
																												--"00110000000000000000000000110011",--59 JMP IMM go to 54



-- 1
"00000100000111100000000000000001",	--49	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--50	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000000001",--51 SHL R10 R13 1
"00011001010011100000000000011111",--52 SHR R10 R14 31
"00000001101011100101000000010000",--53 ADD R13 R14 R10
"00110000000000000000000011101011",	--54	Jmp	��

-- 2
"00000100000111100000000000000010",	--55	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--56	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000000010",--57 SHL R10 R13 2
"00011001010011100000000000011110",--58 SHR R10 R14 30
"00000001101011100101000000010000",--59 ADD R13 R14 R10
"00110000000000000000000011101011",	--60	Jmp	��
--3
"00000100000111100000000000000011",	--61	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--62	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000000011",--63 SHL R10 R13 3
"00011001010011100000000000011101",--64 SHR R10 R14 29
"00000001101011100101000000010000",--65 ADD R13 R14 R10
"00110000000000000000000011101011",	--66	Jmp	��
--4
"00000100000111100000000000000100",	--67	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--68	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000000100",--69 SHL R10 R13 4
"00011001010011100000000000011100",--70 SHR R10 R14 28
"00000001101011100101000000010000",--71 ADD R13 R14 R10
"00110000000000000000000011101011",	--72	Jmp	��

--5
"00000100000111100000000000000101",	--73	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--74	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000000101",--75 SHL R10 R13 5
"00011001010011100000000000011011",--76 SHR R10 R14 27
"00000001101011100101000000010000",--77 ADD R13 R14 R10
"00110000000000000000000011101011",	--78	Jmp	��

--6
"00000100000111100000000000000110",	--79	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--80	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000000110",--81 SHL R10 R13 6
"00011001010011100000000000011010",--82 SHR R10 R14 26
"00000001101011100101000000010000",--83 ADD R13 R14 R10
"00110000000000000000000011101011",	--84	Jmp	��

--7
"00000100000111100000000000000111",	--85	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--86	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000000111",--87 SHL R10 R13 7
"00011001010011100000000000011001",--88 SHR R10 R14 25
"00000001101011100101000000010000",--89 ADD R13 R14 R10
"00110000000000000000000011101011",	--90	Jmp	��

--8
"00000100000111100000000000001000",	--91	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--92	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000001000",--93 SHL R10 R13 8
"00011001010011100000000000011000",--94 SHR R10 R14 24
"00000001101011100101000000010000",--95 ADD R13 R14 R10
"00110000000000000000000011101011",	--96	Jmp	��


--9
"00000100000111100000000000001001",	--97	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--98	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000001001",--99 SHL R10 R13 9
"00011001010011100000000000010111",--100 SHR R10 R14 23
"00000001101011100101000000010000",--101 ADD R13 R14 R10
"00110000000000000000000011101011",	--102	Jmp	��

--10
"00000100000111100000000000001010",	--103	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--104	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000001010",--105 SHL R10 R13 10
"00011001010011100000000000010110",--106 SHR R10 R14 22
"00000001101011100101000000010000",--107 ADD R13 R14 R10
"00110000000000000000000011101011",	--108	Jmp	��

--11
"00000100000111100000000000001011",	--109	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--110	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000001011",--111 SHL R10 R13 11
"00011001010011100000000000010101",--112 SHR R10 R14 21
"00000001101011100101000000010000",--113 ADD R13 R14 R10
"00110000000000000000000011101011",	--114	Jmp	��


--12
"00000100000111100000000000001100",	--115	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--116	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000001100",--117 SHL R10 R13 12
"00011001010011100000000000010100",--118 SHR R10 R14 20
"00000001101011100101000000010000",--119 ADD R13 R14 R10
"00110000000000000000000011101011",	--120	Jmp	��


--13
"00000100000111100000000000001101",	--121	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--122	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000001101",--123 SHL R10 R13 13
"00011001010011100000000000010011",--124 SHR R10 R14 19
"00000001101011100101000000010000",--125 ADD R13 R14 R10
"00110000000000000000000011101011",	--126	Jmp	��


--14
"00000100000111100000000000001110",	--127 Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--128	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000001110",--129 SHL R10 R13 14
"00011001010011100000000000010010",--130 SHR R10 R14 18
"00000001101011100101000000010000",--131 ADD R13 R14 R10
"00110000000000000000000011101011",	--132	Jmp	��

--15
"00000100000111100000000000001111",	--133	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--134	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000001111",--135 SHL R10 R13 15
"00011001010011100000000000010001",--136 SHR R10 R14 17
"00000001101011100101000000010000",--137 ADD R13 R14 R10
"00110000000000000000000011101011",	--138	Jmp	��

--16
"00000100000111100000000000010000",	--139	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--140	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000010000",--141 SHL R10 R13 16
"00011001010011100000000000010000",--142 SHR R10 R14 16
"00000001101011100101000000010000",--143 ADD R13 R14 R10
"00110000000000000000000011101011",	--144	Jmp	��


--17
"00000100000111100000000000010001",	--145	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--146	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000010001",--147 SHL R10 R13 17
"00011001010011100000000000001111",--148 SHR R10 R14 15
"00000001101011100101000000010000",--149 ADD R13 R14 R10
"00110000000000000000000011101011",	--150	Jmp	��

--18
"00000100000111100000000000010010",	--151	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--152	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000010010",--153 SHL R10 R13 18
"00011001010011100000000000001110",--154 SHR R10 R14 14
"00000001101011100101000000010000",--155 ADD R13 R14 R10
"00110000000000000000000011101011",	--156	Jmp	��

--19
"00000100000111100000000000010011",	--157	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--158	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000010011",--159 SHL R10 R13 19
"00011001010011100000000000001101",--160 SHR R10 R14 13
"00000001101011100101000000010000",--161 ADD R13 R14 R10
"00110000000000000000000011101011",	--162	Jmp	��


--20
"00000100000111100000000000010100",	--163	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--164	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000010100",--165 SHL R10 R13 20
"00011001010011100000000000001100",--166 SHR R10 R14 12
"00000001101011100101000000010000",--167 ADD R13 R14 R10
"00110000000000000000000011101011",	--168	Jmp	��

--21
"00000100000111100000000000010101",	--169	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--170	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000010101",--171 SHL R10 R13 21
"00011001010011100000000000001011",--172 SHR R10 R14 11
"00000001101011100101000000010000",--173 ADD R13 R14 R10
"00110000000000000000000011101011",	--174	Jmp	��

--22
"00000100000111100000000000010110",	--175	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--176	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000010110",--177 SHL R10 R13 22
"00011001010011100000000000001010",--178 SHR R10 R14 10
"00000001101011100101000000010000",--179 ADD R13 R14 R10
"00110000000000000000000011101011",	--180	Jmp	��

--23
"00000100000111100000000000010111",	--181	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--182	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000010111",--183 SHL R10 R13 23
"00011001010011100000000000001001",--184 SHR R10 R14 9
"00000001101011100101000000010000",--185 ADD R13 R14 R10
"00110000000000000000000011101011",	--186	Jmp	��

--24
"00000100000111100000000000011000",	--187	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--188	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000011000",--189 SHL R10 R13 24
"00011001010011100000000000001000",--190 SHR R10 R14 8
"00000001101011100101000000010000",--191 ADD R13 R14 R10
"00110000000000000000000011101011",	--192	Jmp	��


--25
"00000100000111100000000000011001",	--193	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--194	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000011001",--195 SHL R10 R13 25
"00011001010011100000000000000111",--196 SHR R10 R14 7
"00000001101011100101000000010000",--197 ADD R13 R14 R10
"00110000000000000000000011101011",	--198	Jmp	��

--26
"00000100000111100000000000011010",	--199	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--200	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000011010",--201 SHL R10 R13 26
"00011001010011100000000000000110",--202 SHR R10 R14 6
"00000001101011100101000000010000",--203 ADD R13 R14 R10
"00110000000000000000000011101011",	--204	Jmp	��


--27
"00000100000111100000000000011011",	--205	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--206	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000011011",--207 SHL R10 R13 27
"00011001010011100000000000000101",--208 SHR R10 R14 5
"00000001101011100101000000010000",--209 ADD R13 R14 R10
"00110000000000000000000011101011",	--210	Jmp	��

--28
"00000100000111100000000000011100",	--211	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--212	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000011100",--213 SHL R10 R13 28
"00011001010011100000000000000100",--214 SHR R10 R14 4
"00000001101011100101000000010000",--215 ADD R13 R14 R10
"00110000000000000000000011101011",	--216	Jmp	��

--29
"00000100000111100000000000011101",	--217	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--218	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000011101",--219 SHL R10 R13 29
"00011001010011100000000000000011",--220 SHR R10 R14 3
"00000001101011100101000000010000",--221 ADD R13 R14 R10
"00110000000000000000000011101011",	--222	Jmp	��

--30
"00000100000111100000000000011110",	--223	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--224	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000011110",--225 SHL R10 R13 30
"00011001010011100000000000000010",--226 SHR R10 R14 2
"00000001101011100101000000010000",--227 ADD R13 R14 R10
"00110000000000000000000011101011",	--228	Jmp	��

--31
"00000100000111100000000000011111",	--229	Addi	0(R00)	counter(R30)		1	
"00101101011111100000000000000100",	--230	Bne	Rotator(R11)	counter(R30)		5	
"00010101010011010000000000011111",--231 SHL R10 R13 31
"00011001010011100000000000000001",--232 SHR R10 R14 1
"00000001101011100101000000010000",--233 ADD R13 R14 R10
"00110000000000000000000011101011",	--234	Jmp	��




"00100000001010100000000000011010",--235 SW R1 R10 IMML branch here  update L[i]
"00000000000010100010100000010000",--236 ADD RO R10 R5
"00000100001000010000000000000001",--237 ADDI R1 R1 1
"00000100010000100000000000000001",--238 ADDI R2 R2 1
"00000100011000110000000000000001",--239 ADDI R3 R3 1
"00101100001101010000000000000001",--240 BNE R1 R21 IMM
"00000000000000000000100000010000",--241 ADD RO RO R1
"00101100010101100000000000000001",--242 BNE R2 R22 IMM
"00000000000000000001000000010000",--243 ADD RO RO R2
"00101000011101110000000000000001",--244 BEQ R3 R22 IMM
"00110000000000000000000000100100",--245 JMP RETURN
"00000000000000000001100000010000",--246 ADD RO RO R3
 


--------------------ENCODE-----------


"00011100000000110000000000000000",	--247	Lw	0(R00)	S[0](R03)		0(Imm��	Load s[0] to R3
"00011100000001000000000000000001",	--248	Lw	0(R00)	S[1](R04)		1(Imm)	Load s[1] to R4
"00000100000001010000000000000000",	--249	Addi	0(R00)	Temp1(R05)		Din(63 downto 48)	
"00010100101001010000000000010000",	--250	Shl	Temp1(R05)	Temp1(R05)		16	Load Din(63 downto 48)
"00000100000001100000000000000000",	--251	Addi	0(R00)	Temp2(R06)		Din(47 downto 32)	
"00010100110001100000000000010000",	--252	Shl	Temp2(R06)	Temp2(R06)		16	
"00011000110001100000000000010000",	--253	Shr	Temp2(R06)	Temp2(R06)		16	Load Din(47 downto 32)
"00000000101001100000100000010000",	--254	Add	Temp1(R05)	Temp2(R06)	A(R01)		Load A
"00000100000001010000000000000000",	--255	Addi	0(R00)	Temp1(R05)		Din(31 downto 16)	
"00010100101001010000000000010000",	--256	Shl	Temp1(R05)	Temp1(R05)		16	Load Din(31 downto 16)
"00000100000001100000000000000000",	--257	Addi	0(R00)	Temp2(R06)		Din(15 downto 0)	
"00010100110001100000000000010000",	--258	Shl	Temp2(R06)	Temp2(R06)		16	
"00011000110001100000000000010000",	--259	Shr	Temp2(R06)	Temp2(R06)		16	Load Din(15 downto 0)
"00000000101001100001000000010000",	--260	Add	Temp1(R05)	Temp2(R06)	B(R02)		Load A


--------------------SELECTION--------------



"00000100000010110000000000000000",	--261	Addi	0(R00)	Mode(R11)			0--encode  1-- decode
"00100100000010110000000110001100",	--262	Blt	0(R00)	Mode(R11)			
"00000000001000110000100000010000",	--263	Add	A(R01)	S[0](R03)	A(R01)		A+s[0]
"00000000010001000001000000010000",	--264	Add	B(R02)	S[1](R04)	B(R02)		B+s[1]
"00000000000000000010100000010000",	--265	Add	0(R00)	0(R00)	I(R05)		Initialize I
"00000100000010100000000000011000",	--266	Addi	0(R00)	24(R10)		24	
"00101000101010100000000110000100",	--267	Beq	I(R05)	24(R10)		388	��
"00000100101001010000000000000010",	--268	Addi	I(R05)	I(R05)		2	I=I+2
"00011100101000110000000000000000",	--269	Lw	I(R05)	S[2*i](R03)		0	Load s[2*i]
"00011100101001000000000000000001",	--270	Lw	I(R05)	S[2*i+1](R04)		1	Load s[2*i+1]
"00000000001000100011000000010010",	--271	And	A(R01)	B(R02)	C(R06)		
"00000000110000000011000000010100",	--272	Nor	C(R06)	0(R00)	C(R06)		
"00000000001000100011100000010011",	--273	Or	A(R01)	B(R02)	D(R07)		
"00000000110001110000100000010010",	--274	And	C(R06)	D(R07)	A(R01)		A Xor B
"00001100010001110000000000011111",	--275	Andi	B(R02)	Rotator(R07)		0000��11111	B(4 downto0)
"00000100000010110000000000000001",	--276	Addi	0(R00)	counter(R11)		1	
"00101100111010110000000000000100",	--277	Bne	Rotator(R07)	counter(R11)		5	
"00010100001010000000000000000001",	--278	Shl	A(R01)	Temp_left(R08)		1	
"00011000001010010000000000011111",	--279	Shr	A(R01)	Temp_right(R09)		31	
"00000001000010010000100000010000",	--280	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--281	Jmp					��
"00000101011010110000000000000001",	--282	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--283	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000000010",	--284	Shl	A(R01)	Temp_left(R08)		2	
"00011000001010010000000000011110",	--285	Shr	A(R01)	Temp_right(R09)		30	
"00000001000010010000100000010000",	--286	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--287	Jmp					��
"00000101011010110000000000000001",	--288	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--289	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000000011",	--290	Shl	A(R01)	Temp_left(R08)		3	
"00011000001010010000000000011101",	--291	Shr	A(R01)	Temp_right(R09)		29	
"00000001000010010000100000010000",	--292	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--293	Jmp					��
"00000101011010110000000000000001",	--294	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--295	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000000100",	--296	Shl	A(R01)	Temp_left(R08)		4	
"00011000001010010000000000011100",	--297	Shr	A(R01)	Temp_right(R09)		28	
"00000001000010010000100000010000",	--298	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--299	Jmp					��
"00000101011010110000000000000001",	--300	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--301	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000000101",	--302	Shl	A(R01)	Temp_left(R08)		5	
"00011000001010010000000000011011",	--303	Shr	A(R01)	Temp_right(R09)		27	
"00000001000010010000100000010000",	--304	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--305	Jmp					��
"00000101011010110000000000000001",	--306	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--307	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000000110",	--308	Shl	A(R01)	Temp_left(R08)		6	
"00011000001010010000000000011010",	--309	Shr	A(R01)	Temp_right(R09)		26	
"00000001000010010000100000010000",	--310	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--311	Jmp					��
"00000101011010110000000000000001",	--312	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--313	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000000111",	--314	Shl	A(R01)	Temp_left(R08)		7	
"00011000001010010000000000011001",	--315	Shr	A(R01)	Temp_right(R09)		25	
"00000001000010010000100000010000",	--316	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--317	Jmp					��
"00000101011010110000000000000001",	--318	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--319	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000001000",	--320	Shl	A(R01)	Temp_left(R08)		8	
"00011000001010010000000000011000",	--321	Shr	A(R01)	Temp_right(R09)		24	
"00000001000010010000100000010000",	--322	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--323	Jmp					��
"00000101011010110000000000000001",	--324	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--325	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000001001",	--326	Shl	A(R01)	Temp_left(R08)		9	
"00011000001010010000000000010111",	--327	Shr	A(R01)	Temp_right(R09)		23	
"00000001000010010000100000010000",	--328	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--329	Jmp					��
"00000101011010110000000000000001",	--330	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--331	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000001010",	--332	Shl	A(R01)	Temp_left(R08)		10	
"00011000001010010000000000010110",	--333	Shr	A(R01)	Temp_right(R09)		22	
"00000001000010010000100000010000",	--334	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--335	Jmp					��
"00000101011010110000000000000001",	--336	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--337	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000001011",	--338	Shl	A(R01)	Temp_left(R08)		11	
"00011000001010010000000000010101",	--339	Shr	A(R01)	Temp_right(R09)		21	
"00000001000010010000100000010000",	--340	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--341	Jmp					��
"00000101011010110000000000000001",	--342	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--343	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000001100",	--344	Shl	A(R01)	Temp_left(R08)		12	
"00011000001010010000000000010100",	--345	Shr	A(R01)	Temp_right(R09)		20	
"00000001000010010000100000010000",	--346	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--347	Jmp					��
"00000101011010110000000000000001",	--348	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--349	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000001101",	--350	Shl	A(R01)	Temp_left(R08)		13	
"00011000001010010000000000010011",	--351	Shr	A(R01)	Temp_right(R09)		19	
"00000001000010010000100000010000",	--352	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--353	Jmp					��
"00000101011010110000000000000001",	--354	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--355	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000001110",	--356	Shl	A(R01)	Temp_left(R08)		14	
"00011000001010010000000000010010",	--357	Shr	A(R01)	Temp_right(R09)		18	
"00000001000010010000100000010000",	--358	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--359	Jmp					��
"00000101011010110000000000000001",	--360	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--361	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000001111",	--362	Shl	A(R01)	Temp_left(R08)		15	
"00011000001010010000000000010001",	--363	Shr	A(R01)	Temp_right(R09)		17	
"00000001000010010000100000010000",	--364	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--365	Jmp					��
"00000101011010110000000000000001",	--366	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--367	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000010000",	--368	Shl	A(R01)	Temp_left(R08)		16	
"00011000001010010000000000010000",	--369	Shr	A(R01)	Temp_right(R09)		16	
"00000001000010010000100000010000",	--370	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--371	Jmp					��
"00000101011010110000000000000001",	--372	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--373	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000010001",	--374	Shl	A(R01)	Temp_left(R08)		17	
"00011000001010010000000000001111",	--375	Shr	A(R01)	Temp_right(R09)		15	
"00000001000010010000100000010000",	--376	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--377	Jmp					��
"00000101011010110000000000000001",	--378	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--379	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000010010",	--380	Shl	A(R01)	Temp_left(R08)		18	
"00011000001010010000000000001110",	--381	Shr	A(R01)	Temp_right(R09)		14	
"00000001000010010000100000010000",	--382	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--383	Jmp					��
"00000101011010110000000000000001",	--384	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--385	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000010011",	--386	Shl	A(R01)	Temp_left(R08)		19	
"00011000001010010000000000001101",	--387	Shr	A(R01)	Temp_right(R09)		13	
"00000001000010010000100000010000",	--388	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--389	Jmp					��
"00000101011010110000000000000001",	--390	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--391	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000010100",	--392	Shl	A(R01)	Temp_left(R08)		20	
"00011000001010010000000000001100",	--393	Shr	A(R01)	Temp_right(R09)		12	
"00000001000010010000100000010000",	--394	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--395	Jmp					��
"00000101011010110000000000000001",	--396	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--397	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000010101",	--398	Shl	A(R01)	Temp_left(R08)		21	
"00011000001010010000000000001011",	--399	Shr	A(R01)	Temp_right(R09)		11	
"00000001000010010000100000010000",	--400	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--401	Jmp					��
"00000101011010110000000000000001",	--402	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--403	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000010110",	--404	Shl	A(R01)	Temp_left(R08)		22	
"00011000001010010000000000001010",	--405	Shr	A(R01)	Temp_right(R09)		10	
"00000001000010010000100000010000",	--406	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--407	Jmp					��
"00000101011010110000000000000001",	--408	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--409	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000010111",	--410	Shl	A(R01)	Temp_left(R08)		23	
"00011000001010010000000000001001",	--411	Shr	A(R01)	Temp_right(R09)		9	
"00000001000010010000100000010000",	--412	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--413	Jmp					��
"00000101011010110000000000000001",	--414	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--415	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000011000",	--416	Shl	A(R01)	Temp_left(R08)		24	
"00011000001010010000000000001000",	--417	Shr	A(R01)	Temp_right(R09)		8	
"00000001000010010000100000010000",	--418	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--419	Jmp					��
"00000101011010110000000000000001",	--420	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--421	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000011001",	--422	Shl	A(R01)	Temp_left(R08)		25	
"00011000001010010000000000000111",	--423	Shr	A(R01)	Temp_right(R09)		7	
"00000001000010010000100000010000",	--424	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--425	Jmp					��
"00000101011010110000000000000001",	--426	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--427	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000011010",	--428	Shl	A(R01)	Temp_left(R08)		26	
"00011000001010010000000000000110",	--429	Shr	A(R01)	Temp_right(R09)		6	
"00000001000010010000100000010000",	--430	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--431	Jmp					��
"00000101011010110000000000000001",	--432	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--433	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000011011",	--434	Shl	A(R01)	Temp_left(R08)		27	
"00011000001010010000000000000101",	--435	Shr	A(R01)	Temp_right(R09)		5	
"00000001000010010000100000010000",	--436	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--437	Jmp					��
"00000101011010110000000000000001",	--438	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--439	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000011100",	--440	Shl	A(R01)	Temp_left(R08)		28	
"00011000001010010000000000000100",	--441	Shr	A(R01)	Temp_right(R09)		4	
"00000001000010010000100000010000",	--442	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--443	Jmp					��
"00000101011010110000000000000001",	--444	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--445	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000011101",	--446	Shl	A(R01)	Temp_left(R08)		29	
"00011000001010010000000000000011",	--447	Shr	A(R01)	Temp_right(R09)		3	
"00000001000010010000100000010000",	--448	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--449	Jmp					��
"00000101011010110000000000000001",	--450	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--451	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000011110",	--452	Shl	A(R01)	Temp_left(R08)		30	
"00011000001010010000000000000010",	--453	Shr	A(R01)	Temp_right(R09)		2	
"00000001000010010000100000010000",	--454	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--455	Jmp					��
"00000101011010110000000000000001",	--456	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--457	Bne	Rotator(R07)	counter(R11)		4	
"00010100001010000000000000011111",	--458	Shl	A(R01)	Temp_left(R08)		31	
"00011000001010010000000000000001",	--459	Shr	A(R01)	Temp_right(R09)		1	
"00000001000010010000100000010000",	--460	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000000111001110",	--461	Jmp					��
"00000000001000110000100000010000",	--462	Add	A(R01)	S[2*i](R03)	A(R01)	��	A=xxx+s[2*i]
"00000000001000100011000000010010",	--463	And	A(R01)	B(R02)	C(R06)		
"00000000110000000011000000010100",	--464	Nor	C(R06)	0(R00)	C(R06)		
"00000000001000100011100000010011",	--465	Or	A(R01)	B(R02)	D(R07)		
"00000000110001110001000000010010",	--466	And	C(R06)	D(R07)	B(R02)		A Xor B
"00001100001001110000000000011111",	--467	Andi	A(R01)	Rotator(R07)		0000��11111	A(4 downto0)
"00000100000010110000000000000001",	--468	Addi	0(R00)	counter(R11)		1	
"00101100111010110000000000000100",	--469	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000000001",	--470	Shl	B(R02)	Temp_left(R08)		1	
"00011000010010010000000000011111",	--471	Shr	B(R02)	Temp_right(R09)		31	
"00000001000010010001000000010000",	--472	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--473	Jmp					��
"00000101011010110000000000000001",	--474	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--475	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000000010",	--476	Shl	B(R02)	Temp_left(R08)		2	
"00011000010010010000000000011110",	--477	Shr	B(R02)	Temp_right(R09)		30	
"00000001000010010001000000010000",	--478	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--479	Jmp					��
"00000101011010110000000000000001",	--480	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--481	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000000011",	--482	Shl	B(R02)	Temp_left(R08)		3	
"00011000010010010000000000011101",	--483	Shr	B(R02)	Temp_right(R09)		29	
"00000001000010010001000000010000",	--484	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--485	Jmp					��
"00000101011010110000000000000001",	--486	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--487	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000000100",	--488	Shl	B(R02)	Temp_left(R08)		4	
"00011000010010010000000000011100",	--489	Shr	B(R02)	Temp_right(R09)		28	
"00000001000010010001000000010000",	--490	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--491	Jmp					��
"00000101011010110000000000000001",	--492	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--493	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000000101",	--494	Shl	B(R02)	Temp_left(R08)		5	
"00011000010010010000000000011011",	--495	Shr	B(R02)	Temp_right(R09)		27	
"00000001000010010001000000010000",	--496	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--497	Jmp					��
"00000101011010110000000000000001",	--498	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--499	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000000110",	--500	Shl	B(R02)	Temp_left(R08)		6	
"00011000010010010000000000011010",	--501	Shr	B(R02)	Temp_right(R09)		26	
"00000001000010010001000000010000",	--502	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--503	Jmp					��
"00000101011010110000000000000001",	--504	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--505	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000000111",	--506	Shl	B(R02)	Temp_left(R08)		7	
"00011000010010010000000000011001",	--507	Shr	B(R02)	Temp_right(R09)		25	
"00000001000010010001000000010000",	--508	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--509	Jmp					��
"00000101011010110000000000000001",	--510	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--511	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000001000",	--512	Shl	B(R02)	Temp_left(R08)		8	
"00011000010010010000000000011000",	--513	Shr	B(R02)	Temp_right(R09)		24	
"00000001000010010001000000010000",	--514	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--515	Jmp					��
"00000101011010110000000000000001",	--516	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--517	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000001001",	--518	Shl	B(R02)	Temp_left(R08)		9	
"00011000010010010000000000010111",	--519	Shr	B(R02)	Temp_right(R09)		23	
"00000001000010010001000000010000",	--520	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--521	Jmp					��
"00000101011010110000000000000001",	--522	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--523	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000001010",	--524	Shl	B(R02)	Temp_left(R08)		10	
"00011000010010010000000000010110",	--525	Shr	B(R02)	Temp_right(R09)		22	
"00000001000010010001000000010000",	--526	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--527	Jmp					��
"00000101011010110000000000000001",	--528	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--529	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000001011",	--530	Shl	B(R02)	Temp_left(R08)		11	
"00011000010010010000000000010101",	--531	Shr	B(R02)	Temp_right(R09)		21	
"00000001000010010001000000010000",	--532	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--533	Jmp					��
"00000101011010110000000000000001",	--534	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--535	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000001100",	--536	Shl	B(R02)	Temp_left(R08)		12	
"00011000010010010000000000010100",	--537	Shr	B(R02)	Temp_right(R09)		20	
"00000001000010010001000000010000",	--538	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--539	Jmp					��
"00000101011010110000000000000001",	--540	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--541	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000001101",	--542	Shl	B(R02)	Temp_left(R08)		13	
"00011000010010010000000000010011",	--543	Shr	B(R02)	Temp_right(R09)		19	
"00000001000010010001000000010000",	--544	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--545	Jmp					��
"00000101011010110000000000000001",	--546	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--547	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000001110",	--548	Shl	B(R02)	Temp_left(R08)		14	
"00011000010010010000000000010010",	--549	Shr	B(R02)	Temp_right(R09)		18	
"00000001000010010001000000010000",	--550	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--551	Jmp					��
"00000101011010110000000000000001",	--552	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--553	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000001111",	--554	Shl	B(R02)	Temp_left(R08)		15	
"00011000010010010000000000010001",	--555	Shr	B(R02)	Temp_right(R09)		17	
"00000001000010010001000000010000",	--556	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--557	Jmp					��
"00000101011010110000000000000001",	--558	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--559	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000010000",	--560	Shl	B(R02)	Temp_left(R08)		16	
"00011000010010010000000000010000",	--561	Shr	B(R02)	Temp_right(R09)		16	
"00000001000010010001000000010000",	--562	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--563	Jmp					��
"00000101011010110000000000000001",	--564	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--565	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000010001",	--566	Shl	B(R02)	Temp_left(R08)		17	
"00011000010010010000000000001111",	--567	Shr	B(R02)	Temp_right(R09)		15	
"00000001000010010001000000010000",	--568	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--569	Jmp					��
"00000101011010110000000000000001",	--570	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--571	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000010010",	--572	Shl	B(R02)	Temp_left(R08)		18	
"00011000010010010000000000001110",	--573	Shr	B(R02)	Temp_right(R09)		14	
"00000001000010010001000000010000",	--574	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--575	Jmp					��
"00000101011010110000000000000001",	--576	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--577	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000010011",	--578	Shl	B(R02)	Temp_left(R08)		19	
"00011000010010010000000000001101",	--579	Shr	B(R02)	Temp_right(R09)		13	
"00000001000010010001000000010000",	--580	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--581	Jmp					��
"00000101011010110000000000000001",	--582	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--583	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000010100",	--584	Shl	B(R02)	Temp_left(R08)		20	
"00011000010010010000000000001100",	--585	Shr	B(R02)	Temp_right(R09)		12	
"00000001000010010001000000010000",	--586	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--587	Jmp					��
"00000101011010110000000000000001",	--588	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--589	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000010101",	--590	Shl	B(R02)	Temp_left(R08)		21	
"00011000010010010000000000001011",	--591	Shr	B(R02)	Temp_right(R09)		11	
"00000001000010010001000000010000",	--592	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--593	Jmp					��
"00000101011010110000000000000001",	--594	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--595	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000010110",	--596	Shl	B(R02)	Temp_left(R08)		22	
"00011000010010010000000000001010",	--597	Shr	B(R02)	Temp_right(R09)		10	
"00000001000010010001000000010000",	--598	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--599	Jmp					��
"00000101011010110000000000000001",	--600	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--601	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000010111",	--602	Shl	B(R02)	Temp_left(R08)		23	
"00011000010010010000000000001001",	--603	Shr	B(R02)	Temp_right(R09)		9	
"00000001000010010001000000010000",	--604	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--605	Jmp					��
"00000101011010110000000000000001",	--606	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--607	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000011000",	--608	Shl	B(R02)	Temp_left(R08)		24	
"00011000010010010000000000001000",	--609	Shr	B(R02)	Temp_right(R09)		8	
"00000001000010010001000000010000",	--610	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--611	Jmp					��
"00000101011010110000000000000001",	--612	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--613	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000011001",	--614	Shl	B(R02)	Temp_left(R08)		25	
"00011000010010010000000000000111",	--615	Shr	B(R02)	Temp_right(R09)		7	
"00000001000010010001000000010000",	--616	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--617	Jmp					��
"00000101011010110000000000000001",	--618	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--619	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000011010",	--620	Shl	B(R02)	Temp_left(R08)		26	
"00011000010010010000000000000110",	--621	Shr	B(R02)	Temp_right(R09)		6	
"00000001000010010001000000010000",	--622	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--623	Jmp					��
"00000101011010110000000000000001",	--624	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--625	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000011011",	--626	Shl	B(R02)	Temp_left(R08)		27	
"00011000010010010000000000000101",	--627	Shr	B(R02)	Temp_right(R09)		5	
"00000001000010010001000000010000",	--628	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--629	Jmp					��
"00000101011010110000000000000001",	--630	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--631	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000011100",	--632	Shl	B(R02)	Temp_left(R08)		28	
"00011000010010010000000000000100",	--633	Shr	B(R02)	Temp_right(R09)		4	
"00000001000010010001000000010000",	--634	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--635	Jmp					��
"00000101011010110000000000000001",	--636	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--637	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000011101",	--638	Shl	B(R02)	Temp_left(R08)		29	
"00011000010010010000000000000011",	--639	Shr	B(R02)	Temp_right(R09)		3	
"00000001000010010001000000010000",	--640	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--641	Jmp					��
"00000101011010110000000000000001",	--642	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--643	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000011110",	--644	Shl	B(R02)	Temp_left(R08)		30	
"00011000010010010000000000000010",	--645	Shr	B(R02)	Temp_right(R09)		2	
"00000001000010010001000000010000",	--646	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--647	Jmp					��
"00000101011010110000000000000001",	--648	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--649	Bne	Rotator(R07)	counter(R11)		4	
"00010100010010000000000000011111",	--650	Shl	B(R02)	Temp_left(R08)		31	
"00011000010010010000000000000001",	--651	Shr	B(R02)	Temp_right(R09)		1	
"00000001000010010001000000010000",	--652	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001010001110",	--653	Jmp					��
"00000000010001000001000000010000",	--654	Add	B(R02)	S[2*i+1](R04)	B(R02)	��	B=xxx+s[2*i+1]
"00110000000000000000000100001011",	--655	Jmp				��	Loop back
"00000000001000001111100000010000",	--656	Add	A(R01)	0(R00)	Dec_out(R31)		
"00000000010000001111000000010000",	--657	Add	B(R02)	0(R00)	Dec_out(R30)		
"11111111111111111111111111111111",	--658	Halt					


------------DECODE---------------------


"00000100000010100000000000011000",	--659	Addi	0(R00)	24(R10)		24	Start of DEC
"00000000000010100010100000010000",	--660	Add	0(R00)	24(R10)	I(R05)		Initialize I
"00101000101000000000000110000100",	--661	Beq	I(R05)	0(R00)		388	��
"00011100101000110000000000000000",	--662	Lw	I(R05)	S[2*i](R03)		0	Load s[2*i]
"00011100101001000000000000000001",	--663	Lw	I(R05)	S[2*i+1](R04)		1	Load s[2*i+1]
"00001000101001010000000000000010",	--664	Subi	I(R05)	I(R05)		2	I=I-2
"00000000010001000001000000010001",	--665	Sub	B(R02)	S[2*i+1](R04)	B(R02)		 B=xxx-s[2*i+1]
"00001100001001110000000000011111",	--666	Andi	A(R01)	Rotator(R07)		0000��11111	A(4 downto0)
"00000100000010110000000000000001",	--667	Addi	0(R00)	counter(R11)		1	
"00101100111010110000000000000100",	--668	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000000001",	--669	Shr	B(R02)	Temp_left(R08)		1	
"00010100010010010000000000011111",	--670	Shl	B(R02)	Temp_right(R09)		31	
"00000001000010010001000000010000",	--671	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--672	Jmp					��
"00000101011010110000000000000001",	--673	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--674	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000000010",	--675	Shr	B(R02)	Temp_left(R08)		2	
"00010100010010010000000000011110",	--676	Shl	B(R02)	Temp_right(R09)		30	
"00000001000010010001000000010000",	--677	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--678	Jmp					��
"00000101011010110000000000000001",	--679	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--680	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000000011",	--681	Shr	B(R02)	Temp_left(R08)		3	
"00010100010010010000000000011101",	--682	Shl	B(R02)	Temp_right(R09)		29	
"00000001000010010001000000010000",	--683	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--684	Jmp					��
"00000101011010110000000000000001",	--685	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--686	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000000100",	--687	Shr	B(R02)	Temp_left(R08)		4	
"00010100010010010000000000011100",	--688	Shl	B(R02)	Temp_right(R09)		28	
"00000001000010010001000000010000",	--689	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--690	Jmp					��
"00000101011010110000000000000001",	--691	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--692	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000000101",	--693	Shr	B(R02)	Temp_left(R08)		5	
"00010100010010010000000000011011",	--694	Shl	B(R02)	Temp_right(R09)		27	
"00000001000010010001000000010000",	--695	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--696	Jmp					��
"00000101011010110000000000000001",	--697	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--698	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000000110",	--699	Shr	B(R02)	Temp_left(R08)		6	
"00010100010010010000000000011010",	--700	Shl	B(R02)	Temp_right(R09)		26	
"00000001000010010001000000010000",	--701	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--702	Jmp					��
"00000101011010110000000000000001",	--703	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--704	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000000111",	--705	Shr	B(R02)	Temp_left(R08)		7	
"00010100010010010000000000011001",	--706	Shl	B(R02)	Temp_right(R09)		25	
"00000001000010010001000000010000",	--707	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--708	Jmp					��
"00000101011010110000000000000001",	--709	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--710	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000001000",	--711	Shr	B(R02)	Temp_left(R08)		8	
"00010100010010010000000000011000",	--712	Shl	B(R02)	Temp_right(R09)		24	
"00000001000010010001000000010000",	--713	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--714	Jmp					��
"00000101011010110000000000000001",	--715	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--716	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000001001",	--717	Shr	B(R02)	Temp_left(R08)		9	
"00010100010010010000000000010111",	--718	Shl	B(R02)	Temp_right(R09)		23	
"00000001000010010001000000010000",	--719	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--720	Jmp					��
"00000101011010110000000000000001",	--721	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--722	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000001010",	--723	Shr	B(R02)	Temp_left(R08)		10	
"00010100010010010000000000010110",	--724	Shl	B(R02)	Temp_right(R09)		22	
"00000001000010010001000000010000",	--725	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--726	Jmp					��
"00000101011010110000000000000001",	--727	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--728	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000001011",	--729	Shr	B(R02)	Temp_left(R08)		11	
"00010100010010010000000000010101",	--730	Shl	B(R02)	Temp_right(R09)		21	
"00000001000010010001000000010000",	--731	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--732	Jmp					��
"00000101011010110000000000000001",	--733	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--734	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000001100",	--735	Shr	B(R02)	Temp_left(R08)		12	
"00010100010010010000000000010100",	--736	Shl	B(R02)	Temp_right(R09)		20	
"00000001000010010001000000010000",	--737	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--738	Jmp					��
"00000101011010110000000000000001",	--739	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--740	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000001101",	--741	Shr	B(R02)	Temp_left(R08)		13	
"00010100010010010000000000010011",	--742	Shl	B(R02)	Temp_right(R09)		19	
"00000001000010010001000000010000",	--743	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--744	Jmp					��
"00000101011010110000000000000001",	--745	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--746	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000001110",	--747	Shr	B(R02)	Temp_left(R08)		14	
"00010100010010010000000000010010",	--748	Shl	B(R02)	Temp_right(R09)		18	
"00000001000010010001000000010000",	--749	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--750	Jmp					��
"00000101011010110000000000000001",	--751	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--752	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000001111",	--753	Shr	B(R02)	Temp_left(R08)		15	
"00010100010010010000000000010001",	--754	Shl	B(R02)	Temp_right(R09)		17	
"00000001000010010001000000010000",	--755	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--756	Jmp					��
"00000101011010110000000000000001",	--757	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--758	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000010000",	--759	Shr	B(R02)	Temp_left(R08)		16	
"00010100010010010000000000010000",	--760	Shl	B(R02)	Temp_right(R09)		16	
"00000001000010010001000000010000",	--761	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--762	Jmp					��
"00000101011010110000000000000001",	--763	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--764	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000010001",	--765	Shr	B(R02)	Temp_left(R08)		17	
"00010100010010010000000000001111",	--766	Shl	B(R02)	Temp_right(R09)		15	
"00000001000010010001000000010000",	--767	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--768	Jmp					��
"00000101011010110000000000000001",	--769	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--770	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000010010",	--771	Shr	B(R02)	Temp_left(R08)		18	
"00010100010010010000000000001110",	--772	Shl	B(R02)	Temp_right(R09)		14	
"00000001000010010001000000010000",	--773	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--774	Jmp					��
"00000101011010110000000000000001",	--775	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--776	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000010011",	--777	Shr	B(R02)	Temp_left(R08)		19	
"00010100010010010000000000001101",	--778	Shl	B(R02)	Temp_right(R09)		13	
"00000001000010010001000000010000",	--779	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--780	Jmp					��
"00000101011010110000000000000001",	--781	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--782	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000010100",	--783	Shr	B(R02)	Temp_left(R08)		20	
"00010100010010010000000000001100",	--784	Shl	B(R02)	Temp_right(R09)		12	
"00000001000010010001000000010000",	--785	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--786	Jmp					��
"00000101011010110000000000000001",	--787	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--788	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000010101",	--789	Shr	B(R02)	Temp_left(R08)		21	
"00010100010010010000000000001011",	--790	Shl	B(R02)	Temp_right(R09)		11	
"00000001000010010001000000010000",	--791	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--792	Jmp					��
"00000101011010110000000000000001",	--793	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--794	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000010110",	--795	Shr	B(R02)	Temp_left(R08)		22	
"00010100010010010000000000001010",	--796	Shl	B(R02)	Temp_right(R09)		10	
"00000001000010010001000000010000",	--797	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--798	Jmp					��
"00000101011010110000000000000001",	--799	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--800	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000010111",	--801	Shr	B(R02)	Temp_left(R08)		23	
"00010100010010010000000000001001",	--802	Shl	B(R02)	Temp_right(R09)		9	
"00000001000010010001000000010000",	--803	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--804	Jmp					��
"00000101011010110000000000000001",	--805	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--806	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000011000",	--807	Shr	B(R02)	Temp_left(R08)		24	
"00010100010010010000000000001000",	--808	Shl	B(R02)	Temp_right(R09)		8	
"00000001000010010001000000010000",	--809	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--810	Jmp					��
"00000101011010110000000000000001",	--811	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--812	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000011001",	--813	Shr	B(R02)	Temp_left(R08)		25	
"00010100010010010000000000000111",	--814	Shl	B(R02)	Temp_right(R09)		7	
"00000001000010010001000000010000",	--815	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--816	Jmp					��
"00000101011010110000000000000001",	--817	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--818	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000011010",	--819	Shr	B(R02)	Temp_left(R08)		26	
"00010100010010010000000000000110",	--820	Shl	B(R02)	Temp_right(R09)		6	
"00000001000010010001000000010000",	--821	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--822	Jmp					��
"00000101011010110000000000000001",	--823	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--824	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000011011",	--825	Shr	B(R02)	Temp_left(R08)		27	
"00010100010010010000000000000101",	--826	Shl	B(R02)	Temp_right(R09)		5	
"00000001000010010001000000010000",	--827	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001101010101",	--828	Jmp					��
"00000101011010110000000000000001",	--829	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--830	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000011100",	--831	Shr	B(R02)	Temp_left(R08)		28	
"00010100010010010000000000000100",	--832	Shl	B(R02)	Temp_right(R09)		4	
"00000001000010010001000000010000",	--833	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--834	Jmp					��
"00000101011010110000000000000001",	--835	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--836	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000011101",	--837	Shr	B(R02)	Temp_left(R08)		29	
"00010100010010010000000000000011",	--838	Shl	B(R02)	Temp_right(R09)		3	
"00000001000010010001000000010000",	--839	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate A
"00110000000000000000001101010101",	--840	Jmp					��
"00000101011010110000000000000001",	--841	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--842	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000011110",	--843	Shr	B(R02)	Temp_left(R08)		30	
"00010100010010010000000000000010",	--844	Shl	B(R02)	Temp_right(R09)		2	
"00000001000010010001000000010000",	--845	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--846	Jmp					��
"00000101011010110000000000000001",	--847	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--848	Bne	Rotator(R07)	counter(R11)		4	
"00011000010010000000000000011111",	--849	Shr	B(R02)	Temp_left(R08)		31	
"00010100010010010000000000000001",	--850	Shl	B(R02)	Temp_right(R09)		1	
"00000001000010010001000000010000",	--851	Add	Temp_left(R08)	Temp_right(R09)	B(R02)		Round rotate B
"00110000000000000000001101010101",	--852	Jmp					��
"00000000001000100011000000010010",	--853	And	A(R01)	B(R02)	C(R06)	��	
"00000000110000000011000000010100",	--854	Nor	C(R06)	0(R00)	C(R06)		
"00000000001000100011100000010011",	--855	Or	A(R01)	B(R02)	D(R07)		
"00000000110001110001000000010010",	--856	And	C(R06)	D(R07)	B(R02)		B = B Xor A
"00000000001000110000100000010001",	--857	Sub	A(R01)	S[2*i](R03)	A(R01)		A=xxx-s[2*i]
"00001100010001110000000000011111",	--858	Andi	B(R02)	Rotator(R07)		0000��11111	B(4 downto0)
"00000100000010110000000000000001",	--859	Addi	0(R00)	counter(R11)		1	
"00101100111010110000000000000100",	--860	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000000001",	--861	Shr	A(R01)	Temp_left(R08)		1	
"00010100001010010000000000011111",	--862	Shl	A(R01)	Temp_right(R09)		31	
"00000001000010010000100000010000",	--863	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--864	Jmp					��
"00000101011010110000000000000001",	--865	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--866	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000000010",	--867	Shr	A(R01)	Temp_left(R08)		2	
"00010100001010010000000000011110",	--868	Shl	A(R01)	Temp_right(R09)		30	
"00000001000010010000100000010000",	--869	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--870	Jmp					��
"00000101011010110000000000000001",	--871	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--872	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000000011",	--873	Shr	A(R01)	Temp_left(R08)		3	
"00010100001010010000000000011101",	--874	Shl	A(R01)	Temp_right(R09)		29	
"00000001000010010000100000010000",	--875	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--876	Jmp					��
"00000101011010110000000000000001",	--877	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--878	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000000100",	--879	Shr	A(R01)	Temp_left(R08)		4	
"00010100001010010000000000011100",	--880	Shl	A(R01)	Temp_right(R09)		28	
"00000001000010010000100000010000",	--881	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--882	Jmp					��
"00000101011010110000000000000001",	--883	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--884	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000000101",	--885	Shr	A(R01)	Temp_left(R08)		5	
"00010100001010010000000000011011",	--886	Shl	A(R01)	Temp_right(R09)		27	
"00000001000010010000100000010000",	--887	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--888	Jmp					��
"00000101011010110000000000000001",	--889	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--890	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000000110",	--891	Shr	A(R01)	Temp_left(R08)		6	
"00010100001010010000000000011010",	--892	Shl	A(R01)	Temp_right(R09)		26	
"00000001000010010000100000010000",	--893	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--894	Jmp					��
"00000101011010110000000000000001",	--895	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--896	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000000111",	--897	Shr	A(R01)	Temp_left(R08)		7	
"00010100001010010000000000011001",	--898	Shl	A(R01)	Temp_right(R09)		25	
"00000001000010010000100000010000",	--899	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--900	Jmp					��
"00000101011010110000000000000001",	--901	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--902	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000001000",	--903	Shr	A(R01)	Temp_left(R08)		8	
"00010100001010010000000000011000",	--904	Shl	A(R01)	Temp_right(R09)		24	
"00000001000010010000100000010000",	--905	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--906	Jmp					��
"00000101011010110000000000000001",	--907	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--908	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000001001",	--909	Shr	A(R01)	Temp_left(R08)		9	
"00010100001010010000000000010111",	--910	Shl	A(R01)	Temp_right(R09)		23	
"00000001000010010000100000010000",	--911	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--912	Jmp					��
"00000101011010110000000000000001",	--913	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--914	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000001010",	--915	Shr	A(R01)	Temp_left(R08)		10	
"00010100001010010000000000010110",	--916	Shl	A(R01)	Temp_right(R09)		22	
"00000001000010010000100000010000",	--917	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--918	Jmp					��
"00000101011010110000000000000001",	--919	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--920	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000001011",	--921	Shr	A(R01)	Temp_left(R08)		11	
"00010100001010010000000000010101",	--922	Shl	A(R01)	Temp_right(R09)		21	
"00000001000010010000100000010000",	--923	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--924	Jmp					��
"00000101011010110000000000000001",	--925	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--926	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000001100",	--927	Shr	A(R01)	Temp_left(R08)		12	
"00010100001010010000000000010100",	--928	Shl	A(R01)	Temp_right(R09)		20	
"00000001000010010000100000010000",	--929	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--930	Jmp					��
"00000101011010110000000000000001",	--931	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--932	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000001101",	--933	Shr	A(R01)	Temp_left(R08)		13	
"00010100001010010000000000010011",	--934	Shl	A(R01)	Temp_right(R09)		19	
"00000001000010010000100000010000",	--935	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--936	Jmp					��
"00000101011010110000000000000001",	--937	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--938	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000001110",	--939	Shr	A(R01)	Temp_left(R08)		14	
"00010100001010010000000000010010",	--940	Shl	A(R01)	Temp_right(R09)		18	
"00000001000010010000100000010000",	--941	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--942	Jmp					��
"00000101011010110000000000000001",	--943	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--944	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000001111",	--945	Shr	A(R01)	Temp_left(R08)		15	
"00010100001010010000000000010001",	--946	Shl	A(R01)	Temp_right(R09)		17	
"00000001000010010000100000010000",	--947	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--948	Jmp					��
"00000101011010110000000000000001",	--949	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--950	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000010000",	--951	Shr	A(R01)	Temp_left(R08)		16	
"00010100001010010000000000010000",	--952	Shl	A(R01)	Temp_right(R09)		16	
"00000001000010010000100000010000",	--953	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--954	Jmp					��
"00000101011010110000000000000001",	--955	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--956	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000010001",	--957	Shr	A(R01)	Temp_left(R08)		17	
"00010100001010010000000000001111",	--958	Shl	A(R01)	Temp_right(R09)		15	
"00000001000010010000100000010000",	--959	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--960	Jmp					��
"00000101011010110000000000000001",	--961	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--962	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000010010",	--963	Shr	A(R01)	Temp_left(R08)		18	
"00010100001010010000000000001110",	--964	Shl	A(R01)	Temp_right(R09)		14	
"00000001000010010000100000010000",	--965	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--966	Jmp					��
"00000101011010110000000000000001",	--967	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--968	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000010011",	--969	Shr	A(R01)	Temp_left(R08)		19	
"00010100001010010000000000001101",	--970	Shl	A(R01)	Temp_right(R09)		13	
"00000001000010010000100000010000",	--971	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--972	Jmp					��
"00000101011010110000000000000001",	--973	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--974	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000010100",	--975	Shr	A(R01)	Temp_left(R08)		20	
"00010100001010010000000000001100",	--976	Shl	A(R01)	Temp_right(R09)		12	
"00000001000010010000100000010000",	--977	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--978	Jmp					��
"00000101011010110000000000000001",	--979	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--980	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000010101",	--981	Shr	A(R01)	Temp_left(R08)		21	
"00010100001010010000000000001011",	--982	Shl	A(R01)	Temp_right(R09)		11	
"00000001000010010000100000010000",	--983	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--984	Jmp					��
"00000101011010110000000000000001",	--985	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--986	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000010110",	--987	Shr	A(R01)	Temp_left(R08)		22	
"00010100001010010000000000001010",	--988	Shl	A(R01)	Temp_right(R09)		10	
"00000001000010010000100000010000",	--989	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--990	Jmp					��
"00000101011010110000000000000001",	--991	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--992	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000010111",	--993	Shr	A(R01)	Temp_left(R08)		23	
"00010100001010010000000000001001",	--994	Shl	A(R01)	Temp_right(R09)		9	
"00000001000010010000100000010000",	--995	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--996	Jmp					��
"00000101011010110000000000000001",	--997	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--998	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000011000",	--999	Shr	A(R01)	Temp_left(R08)		24	
"00010100001010010000000000001000",	--1000	Shl	A(R01)	Temp_right(R09)		8	
"00000001000010010000100000010000",	--1001	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--1002	Jmp					��
"00000101011010110000000000000001",	--1003	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--1004	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000011001",	--1005	Shr	A(R01)	Temp_left(R08)		25	
"00010100001010010000000000000111",	--1006	Shl	A(R01)	Temp_right(R09)		7	
"00000001000010010000100000010000",	--1007	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--1008	Jmp					��
"00000101011010110000000000000001",	--1009	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--1010	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000011010",	--1011	Shr	A(R01)	Temp_left(R08)		26	
"00010100001010010000000000000110",	--1012	Shl	A(R01)	Temp_right(R09)		6	
"00000001000010010000100000010000",	--1013	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--1014	Jmp					��
"00000101011010110000000000000001",	--1015	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--1016	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000011011",	--1017	Shr	A(R01)	Temp_left(R08)		27	
"00010100001010010000000000000101",	--1018	Shl	A(R01)	Temp_right(R09)		5	
"00000001000010010000100000010000",	--1019	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--1020	Jmp					00000000000000010000010101
"00000101011010110000000000000001",	--1021	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--1022	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000011100",	--1023	Shr	A(R01)	Temp_left(R08)		28	
"00010100001010010000000000000100",	--1024	Shl	A(R01)	Temp_right(R09)		4	
"00000001000010010000100000010000",	--1025	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--1026	Jmp					��
"00000101011010110000000000000001",	--1027	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--1028	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000011101",	--1029	Shr	A(R01)	Temp_left(R08)		29	
"00010100001010010000000000000011",	--1030	Shl	A(R01)	Temp_right(R09)		3	
"00000001000010010000100000010000",	--1031	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--1032	Jmp					��
"00000101011010110000000000000001",	--1033	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--1034	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000011110",	--1035	Shr	A(R01)	Temp_left(R08)		30	
"00010100001010010000000000000010",	--1036	Shl	A(R01)	Temp_right(R09)		2	
"00000001000010010000100000010000",	--1037	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--1038	Jmp					��
"00000101011010110000000000000001",	--1039	Addi	counter(R11)	counter(R11)		1	
"00101100111010110000000000000100",	--1040	Bne	Rotator(R07)	counter(R11)		4	
"00011000001010000000000000011111",	--1041	Shr	A(R01)	Temp_left(R08)		31	
"00010100001010010000000000000001",	--1042	Shl	A(R01)	Temp_right(R09)		1	
"00000001000010010000100000010000",	--1043	Add	Temp_left(R08)	Temp_right(R09)	A(R01)		Round rotate A
"00110000000000000000010000010101",	--1044	Jmp					��
"00000000001000100011000000010010",	--1045	And	A(R01)	B(R02)	C(R06)	��	
"00000000110000000011000000010100",	--1046	Nor	C(R06)	0(R00)	C(R06)		
"00000000001000100011100000010011",	--1047	Or	A(R01)	B(R02)	D(R07)		
"00000000110001110000100000010010",	--1048	And	C(R06)	D(R07)	A(R01)		A = A Xor B
"00110000000000000000001010010101",	--1049	Jmp				��	Outer Loop back
"00011100101000110000000000000000",	--1050	Lw	I(R05)	S[0](R03)		0	Load s[0]
"00011100101001000000000000000001",	--1051	Lw	I(R05)	S[1](R04)		1	Load s[1]
"00000000001000110000100000010001",	--1052	Sub	A(R01)	S[0](R03)	A(R01)		A=A-s[0]
"00000000010001000001000000010001",	--1053	Sub	B(R02)	S[1](R04)	B(R02)		 B=B-s[1]
"00000000001000001110100000010000",	--1054	Add	A(R01)	0(R00)	Dec_out(R29)		
"00000000010000001110000000010000",	--1055	Add	B(R02)	0(R00)	Dec_out(R28)		
"11111111111111111111111111111111"	--1056	Halt					
              
 );
 


begin
    imem(3)<="0000010000011110"&skey(31 downto 16);
	 imem(5)<="0000010000011101"&skey(15 downto 0);
	 imem(10)<="0000010000011110"&skey(63 downto 48);
	 imem(12)<="0000010000011101"&skey(47 downto 32);
	 imem(17)<="0000010000011110"&skey(95 downto 80);
	 imem(19)<="0000010000011101"&skey(79 downto 64);
	 imem(24)<="0000010000011110"&skey(127 downto 112);
	 imem(26)<="0000010000011101"&skey(111 downto 96);

	 imem(249)<="0000010000000101"&din(63 downto 48);    --249    Addi    0(R00)    Temp1(R05)        Din(63 downto 48)  
	 imem(251)<="0000010000000110"&din(47 downto 32);    --251    Addi    0(R00)    Temp2(R06)        Din(47 downto 32) 
	 imem(255)<="0000010000000101"&din(31 downto 16);    --255    Addi    0(R00)    Temp1(R05)        Din(31 downto 16)   
	 imem(257)<="0000010000000110"&din(15 downto 0);    --257    Addi    0(R00)    Temp2(R06)        Din(15 downto 0)   
	 
	 imem(261)<="0000010000001011"&"000000000000000"&mode;    --261   Addi    0(R00)    Mode(R11)        Mode  0 for enc; 1 for dec; 
	 		 
    Instruction<=imem(conv_integer(address));
    ins_num <= conv_integer(address);
end Behavioral;