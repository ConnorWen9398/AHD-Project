--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   12:50:51 11/27/2017
-- Design Name:   
-- Module Name:   H:/AVH/dmem/dmem_tb.vhd
-- Project Name:  dmem
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: dmem
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY dmem_tb IS
END dmem_tb;
 
ARCHITECTURE behavior OF dmem_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT dmem
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         address : IN  std_logic_vector(31 downto 0);
         wrtdata : IN  std_logic_vector(31 downto 0);
         wrtmemen : IN  std_logic;
         rddata : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';
   signal address : std_logic_vector(31 downto 0) := (others => '0');
   signal wrtdata : std_logic_vector(31 downto 0) := (others => '0');
   signal wrtmemen : std_logic := '0';

 	--Outputs
   signal rddata : std_logic_vector(31 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: dmem PORT MAP (
          clk => clk,
          reset => reset,
          address => address,
          wrtdata => wrtdata,
          wrtmemen => wrtmemen,
          rddata => rddata
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
      reset<='1';
		address<=x"00000001";
		wrtdata<=x"11111111";
		wrtmemen<='1';
		wait for clk_period;
		reset<='0';
		wrtmemen<='0';
		wait for clk_period;
		wrtmemen<='1';
		wait for clk_period;
		wrtmemen<='0';
		address<=x"00000000";
		wait for clk_period;
		address<=x"00000001";
      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
