
----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:31:53 11/28/2017 
-- Design Name: 
-- Module Name:    InstructionMemory - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity InstructionMemory is
port(
     skey: in std_logic_vector(127 downto 0);
	  din: in std_logic_vector(63 downto 0);
     address: in std_logic_vector(31 downto 0);
	  Instruction: out std_logic_vector(31 downto 0));
	  
end InstructionMemory;

architecture Behavioral of InstructionMemory is

type ramtype3 is array(0 to 160)of std_logic_vector(31 downto 0);
signal imem: ramtype3:=
(
"00000000000000000000100000010000",--0 ADD RO,RO, R1 R1=0
"00000000000000000001000000010000",--1 ADD R0,RO, R2 R2=0
"00000000000000000001100000010000",--2 ADD RO,RO, R3 R3=0
"00000100000111100000000000000000",--3 ****ADDI,RO,R30,skey(31 downto 16) R30=XXX..skey(31 downto 16)
"00010111110111100000000000010000",--4 SHL R30 R30 16 R30=skey(31 downto 16)...000
"00000100000111010000000000000000",--5 ****ADDI,RO,R29,SKEY(15 downto 0) R29=XXX��..skey(15 downto 0)
"00010111101111010000000000010000",--6 SHL R29 R29 16 R29=skey(15 downto 0)��000     remove sign extension
"00011011101111010000000000010000",--7 SHR R29 R29 16 R29=000��..skey(15 downto 0)     remove sign extension
"00000011110111011111000000010000",--8 ADD,R30 R29,R30 R30=skey(31 downto 0) 
"00100000000111100000000000011010",--9 SW RO, R30 offset M[0+offset1]<-R30
"00000100000111100000000000000000",--10 *****ADDI,RO,R30,skey(63 downto 48) R30=XXX..skey(63 downto 48)
"00010111110111100000000000010000",--11 SHL R30 R30 16 R30=skey(63 downto 48)...000
"00000100000111010000000000000000",--12 **** ADDI,RO,R29,SKEY(47 downto 32) R29=XXX��..skey(47 downto 32)
"00010111101111010000000000010000",--13 SHL R29 R29 16 R29=skey(47 downto 32)��000     remove sign extension
"00011011101111010000000000010000",--14 SHR R29 R29 16 R29=000��..skey(47 downto 32)     remove sign extension
"00000011110111011111000000010000",--15 ADD,R30 R29,R30 R30=skey(63 downto 32) 
"00100000000111100000000000011011",--16 SW RO, R30 offset M[0+offset2]<-R30
"00000100000111100000000000000000",--17 ****ADDI,RO,R30,skey(95 downto 80) R30=XXX..skey(95 downto 80)
"00010111110111100000000000010000",--18 SHL R30 R30 16 R30=skey(95 downto 80)...000
"00000100000111010000000000000000",--19 **** ADDI,RO,R29,SKEY(79 downto 64) R29=XXX��..skey(79 downto 64)
"00010111101111010000000000010000",--20 SHL R29 R29 16 R29=skey(79 downto 64)��000     remove sign extension
"00011011101111010000000000010000",--21 SHR R29 R29 16 R29=000��..skey(79 downto 64)     remove sign extension
"00000011110111011111000000010000",--22 ADD,R30 R29,R30 R30=skey(95 downto 64) 
"00100000000111100000000000011100",--23 SW RO, R30 offset M[0+offset3]<-R30
"00000100000111100000000000000000",--24 ******ADDI,RO,R30,skey(127 downto 112) R30=XXX..skey(127 downto 112)
"00010111110111100000000000010000",--25 SHL R30 R30 16 R30=skey(127 downto 112)...000
"00000100000111010000000000000000",--26******* ADDI,RO,R29,SKEY(111 downto 96) R29=XXX��..skey(111 downto 96)
"00010111101111010000000000010000",--27 SHL R29 R29 16 R29=skey(111 downto 96)��000     remove sign extension
"00011011101111010000000000010000",--28 SHR R29 R29 16 R29=000��..skey(111 downto 96)     remove sign extension
"00000011110111011111000000010000",--29 ADD,R30 R29,R30 R30=skey(127 downto 96) 
"00100000000111100000000000011101",--30 SW RO, R30 offset M[0+offset4]<-R30
"00000100000101010000000000000100",--31 ADDI,RO,R21,4 R21=4
"00000100000101100000000000011010",--32 ADDI RO R22,26 R22=26
"00000100000101110000000001001110",--33 ADDI R0 R23,78 R23=78
"00000000000000000010000000010000",--34 ADD RO RO R4 R4=0
"00000000000000000010100000010000",--35 ADD RO RO R5 R5=0
"00011100010010000000000000000000",--36 R8<-MEM[R2+IMM_S) S[i]
"00011100001010010000000000011010",--37 R9<-MEM(R1+IMM_l) L[j]
"00000000100001010011000000010000",--38 ADD R4 R5,R6  A+B
"00000001000001100101000000010000",--39 ADD R8 R6 R10 A+B+S[i]
"00000100000010110000000000000011",--40 ADDI RO R11 3 
"00000000000000000110000000010000",--41 ADD RO RO R12
"00101001011011000000000000000101",--42 BEQ R11 R12 IMM go to 48
"00010101010011010000000000000001",--43 SHL R10 R13 1
"00011001010011100000000000011111",--44 SHR R10 R14 1
"00000001101011100101000000010000",--45 ADD R13 R14 R10  rotate 1 bit of R10, do it 3 times 
"00000101100011000000000000000001",--46 ADDI R12 R12 1
"00110000000000000000000000101010",--47 JMP IMM go to 42
"00100000010010100000000000000000",--48 SW R2 R10 IMM_S branch here update S[i]
"00000000000010100010000000010000",--49 add RO R10 R4 put value of A into R4
"00000000100001010011000000010000",--50 add R4 R5 R6 A + B
"00000001001001100101000000010000",--51 add R9 R6 R10 R10 = L[i] + A + B
"00001100110010110000000000011111",--52 ANDI R6 R11 00....11111
"00000000000000000110000000010000",--53 AND RO RO R12
"00101001011011000000000000000101",--54 bEQ R11 R12 IMM
"00010101010011010000000000000001",--55 SHL R10 R13 1
"00011001010011100000000000011111",--56 SHR R10 R14 31
"00000001101011100101000000010000",--57 ADD R13 R14 R10
"00000101100011000000000000000001",--58 ADDI R12 R12 1
"00110000000000000000000000110110",--59 JMP IMM go to 54
"00100000001010100000000000011010",--60 SW R1 R10 IMML branch here  update L[i]
"00000000000010100010100000010000",--61 ADD RO R10 R5
"00000100001000010000000000000001",--62 ADDI R1 R1 1
"00000100010000100000000000000001",--63 ADDI R2 R2 1
"00000100011000110000000000000001",--64 ADDI R3 R3 1
"00101100001101010000000000000001",--65 BNE R1 R21 IMM
"00000000000000000000100000010000",--66 ADD RO RO R1
"00101100010101100000000000000001",--67 BNE R2 R22 IMM
"00000000000000000001000000010000",--68 ADD RO RO R2
"00101000011101110000000000000001",--69 BEQ R3 R22 IMM
"00110000000000000000000000100100",--70 JMP RETURN
"00000000000000000001100000010000",--71 ADD RO RO R3

----ENCode-----
"00011100000000110000000000000000",    --72    Lw    0(R00)    S[0](R03)        0(Imm��    Load s[0] to R3
"00011100000001000000000000000001",    --73    Lw    0(R00)    S[1](R04)        1(Imm)    Load s[1] to R4
"00000100000001010000000000000000",    --74    Addi    0(R00)    Temp1(R05)        Din(63 downto 48)    
"00010100101001010000000000010000",    --75    Shl    Temp1(R05)    Temp1(R05)        16    Load Din(63 downto 48)
"00000100000001100000000000000000",    --76    Addi    0(R00)    Temp2(R06)        Din(47 downto 32)    
"00010100110001100000000000010000",    --77    Shl    Temp2(R06)    Temp2(R06)        16    
"00011000110001100000000000010000",    --78    Shr    Temp2(R06)    Temp2(R06)        16    Load Din(47 downto 32)
"00000000101001100000100000010000",    --79    Add    Temp1(R05)    Temp2(R06)    A(R01)        Load A
"00000100000001010000000000000000",    --80    Addi    0(R00)    Temp1(R05)        Din(31 downto 16)    
"00010100101001010000000000010000",    --81    Shl    Temp1(R05)    Temp1(R05)        16    Load Din(31 downto 16)
"00000100000001100000000000000000",    --82    Addi    0(R00)    Temp2(R06)        Din(15 downto 0)    
"00010100110001100000000000010000",    --83    Shl    Temp2(R06)    Temp2(R06)        16    
"00011000110001100000000000010000",    --84    Shr    Temp2(R06)    Temp2(R06)        16    Load Din(15 downto 0)
"00000000101001100001000000010000",    --85    Add    Temp1(R05)    Temp2(R06)    B(R02)        Load A
"00000000001000110000100000010000",    --86    Add    A(R01)    S[0](R03)    A(R01)        A+s[0]
"00000000010001000001000000010000",    --87    Add    B(R02)    S[1](R04)    B(R02)        B+s[1]
"00000000000000000010100000010000",    --88    Add    0(R00)    0(R00)    I(R05)        Initialize I
"00000100000010100000000000011000",    --89    Addi    0(R00)    24(R10)        24    
"00101000101010100000000000011100",    --90    Beq    I(R05)    24(R10)        28    ��
"00000100101001010000000000000010",    --91    Addi    I(R05)    I(R05)        2    I=I+2
"00011100101000110000000000000000",    --92    Lw    I(R05)    S[2*i](R03)        0    Load s[2*i]
"00011100101001000000000000000001",    --93    Lw    I(R05)    S[2*i+1](R04)        1    Load s[2*i+1]
"00000000001000100011000000010010",    --94    And    A(R01)    B(R02)    C(R06)        
"00000000110000000011000000010100",    --95    Nor    C(R06)    0(R00)    C(R06)        
"00000000001000100011100000010011",    --96    Or    A(R01)    B(R02)    D(R07)        
"00000000110001110000100000010010",    --97    And    C(R06)    D(R07)    A(R01)        A Xor B
"00001100010001110000000000011111",    --98    Andi    B(R02)    Rotator(R07)        0000��11111    B(4 downto0)
"00101000111000000000000000000101",    --99    Beq    Rotator(R07)    0(R00)        5    ��
"00010100001010000000000000000001",    --100    Shl    A(R01)    Temp_left(R08)        1    
"00011000001010010000000000011111",    --101    Shr    A(R01)    Temp_right(R09)        31    
"00000001000010010000100000010000",    --102    Add    Temp_left(R08)    Temp_right(R09)    A(R01)        Round rotate A
"00001000111001110000000000000001",    --103    Subi    Rotator(R07)    Rotator(R07)        1    
"00110000000000000000000001100011",    --104    Jmp                ��    Loop back
"00000000001000110000100000010000",    --105    Add    A(R01)    S[2*i](R03)    A(R01)        A=xxx+s[2*i]
"00000000001000100011000000010010",    --106    And    A(R01)    B(R02)    C(R06)        
"00000000110000000011000000010100",    --107    Nor    C(R06)    0(R00)    C(R06)        
"00000000001000100011100000010011",    --108    Or    A(R01)    B(R02)    D(R07)        
"00000000110001110001000000010010",    --109    And    C(R06)    D(R07)    B(R02)        A Xor B
"00001100001001110000000000011111",    --110    Andi    A(R01)    Rotator(R07)        0000��11111    A(4 downto0)
"00101000111000000000000000000101",    --111    Beq    Rotator(R07)    0(R00)        5    ��
"00010100010010000000000000000001",    --112    SHL    B(R02)    Temp_left(R08)        1    
"00011000010010010000000000011111",    --113    SHR    B(R02)    Temp_right(R09)        31    
"00000001000010010001000000010000",    --114    Add    Temp_left(R08)    Temp_right(R09)    B(R02)        Round rotate B
"00001000111001110000000000000001",    --115    Subi    Rotator(R07)    Rotator(R07)        1    
"00110000000000000000000001101111",    --116    Jmp                ��    Loop back
"00000000010001000001000000010000",    --117    Add    B(R02)    S[2*i+1](R04)    B(R02)        B=xxx+s[2*i+1]
"00110000000000000000000001011010",    --118    Jmp                ��    Loop back
"00000000001000001111100000010000",	   --119	Add	A(R01)	0(R00)	Dec_out(R31)		
"00000000010000001111000000010000",	   --120	Add	B(R02)	0(R00)	Dec_out(R30)
"00000000000000000010100000010000",    --121    Add    0(R00)    0(R00)    Temp1(R05)        Clear R05
"00000000000000000011000000010000",    --122    Add    0(R00)    0(R00)    Temp1(R06)        Clear R06
"00000100000010100000000000011000",    --123    Addi    0(R00)    24(R10)        24    
"00000000000010100010100000010000",     --124    Add    0(R00)    24(R10)    I(R05)        Initialize I
"00101000101000000000000000011100",     --125    Beq    I(R05)    0(R00)        28    ��
"00011100101000110000000000000000",    --126    Lw    I(R05)    S[2*i](R03)        0    Load s[2*i]
"00011100101001000000000000000001",    --127    Lw    I(R05)    S[2*i+1](R04)        1    Load s[2*i+1]
"00001000101001010000000000000010",    --128    Subi    I(R05)    I(R05)        2    I=I-2
"00000000010001000001000000010001",    --129    Sub    B(R02)    S[2*i+1](R04)    B(R02)        B=xxx-s[2*i+1]
"00001100001001110000000000011111",    --130    Andi    A(R01)    Rotator(R07)        0000��11111    A(4 downto0)
"00101000111000000000000000000101",    --131    Beq    Rotator(R07)    0(R00)        5    ��
"00011000010010000000000000000001",    --132    Shr    B(R02)    Temp_right(R08)        1    
"00010100010010010000000000011111",    --133    Shl    B(R02)    Temp_left(R09)        31    
"00000001000010010001000000010000",    --134    Add    Temp_left(R08)    Temp_right(R09)    B(R02)        Round right rotate B
"00001000111001110000000000000001",    --135    Subi    Rotator(R07)    Rotator(R07)        1    
"00110000000000000000000010000011",    --136    Jmp                ��    Rotate loop1 back
"00000000001000100011000000010010",    --137    And    A(R01)    B(R02)    C(R06)        
"00000000110000000011000000010100",    --138    Nor    C(R06)    0(R00)    C(R06)        
"00000000001000100011100000010011",    --139    Or    A(R01)    B(R02)    D(R07)        
"00000000110001110001000000010010",    --140    And    C(R06)    D(R07)    B(R02)        B= B Xor A
"00000000001000110000100000010001",    --141    Sub    A(R01)    S[2*i](R03)    A(R01)        A=xxx-s[2*i]
"00001100010001110000000000011111",    --142    Andi    B(R02)    Rotator(R07)        0000��11111    B(4 downto0)
"00101000111000000000000000000101",    --143    Beq    Rotator(R07)    0(R00)        5    ��
"00011000001010000000000000000001",    --144    Shr    A(R01)    Temp_right(R08)        1    
"00010100001010010000000000011111",    --145    Shl    A(R01)    Temp_left(R09)        31    
"00000001000010010000100000010000",    --146    Add    Temp_left(R08)    Temp_right(R09)    A(R01)        Round right rotate A
"00001000111001110000000000000001",    --147    Subi    Rotator(R07)    Rotator(R07)        1    
"00110000000000000000000010001111",    --148    Jmp                ��    Rotate loop2 back
"00000000001000100011000000010010",    --149    And    A(R01)    B(R02)    C(R06)        
"00000000110000000011000000010100",    --150    Nor    C(R06)    0(R00)    C(R06)        
"00000000001000100011100000010011",    --151    Or    A(R01)    B(R02)    D(R07)        
"00000000110001110000100000010010",    --152    And    C(R06)    D(R07)    A(R01)        A =A Xor B
"00110000000000000000000001111101",    --153    Jmp                ��    Outer loop back
"00011100000000110000000000000000",    --154    Lw    0(R00)    S[0](R03)        0(Imm��    Load s[0] to R3
"00011100000001000000000000000001",    --155    Lw    0(R00)    S[1](R04)        1(Imm)    Load s[1] to R4
"00000000001000110000100000010001",    --156    Sub    A(R01)    S[0](R03)    A(R01)        A= A - s[0]
"00000000010001000001000000010001",    --157    Sub    B(R02)    S[1](R04)    B(R02)        B= B - s[1]
"00000000001000001110100000010000",    --158    Add    A(R01)    0(R00)    Dec_out(R29)
"00000000010000001110000000010000",    --159    Add    B(R02)    0(R00)    Dec_out(R28)
"11111111111111111111111111111111"      --160   Hal                
 );
signal ins_num : integer;
begin
    imem(3)<="0000010000011110"&skey(31 downto 16);
	 imem(5)<="0000010000011101"&skey(15 downto 0);
	 imem(10)<="0000010000011110"&skey(63 downto 48);
	 imem(12)<="0000010000011101"&skey(47 downto 32);
	 imem(17)<="0000010000011110"&skey(95 downto 80);
	 imem(19)<="0000010000011101"&skey(79 downto 64);
	 imem(24)<="0000010000011110"&skey(127 downto 112);
	 imem(26)<="0000010000011101"&skey(111 downto 96);

	 imem(74)<="0000010000000101"&din(63 downto 48);    --74    Addi    0(R00)    Temp1(R05)        Din(63 downto 48)  
	 imem(76)<="0000010000000110"&din(47 downto 32);    --76    Addi    0(R00)    Temp2(R06)        Din(47 downto 32) 
	 imem(80)<="0000010000000101"&din(31 downto 16);    --80    Addi    0(R00)    Temp1(R05)        Din(31 downto 16)   
	 imem(82)<="0000010000000110"&din(15 downto 0);    --82    Addi    0(R00)    Temp2(R06)        Din(15 downto 0)   
	 		 
    Instruction<=imem(conv_integer(address));
    ins_num <= conv_integer(address);
end Behavioral;